`timescale 1ns/1ns // ????????1ns????????1ns

module flow_led_tb(); // ????

//parameter define
parameter T = 20; // ?????20ns

//reg define
reg sys_clk; // ????
reg sys_rst_n; // ????

//wire define
wire [3:0] led;



//????????
initial begin
sys_clk = 1'b0;
sys_rst_n = 1'b0; // ??
#(T+1) sys_rst_n = 1'b1; // ??21ns???????????
end

//50Mhz????????1/50Mhz=20ns,???10ns???????
always #(T/2) sys_clk = ~sys_clk;

//??flow_led??
flow_led u0_flow_led (
   .sys_clk (sys_clk ),
   .sys_rst_n (sys_rst_n),
   .led (led )
);

endmodule




